library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity sincos_lut_14 is
	port (
		clk_i  : in std_logic;
		addr_i : in std_logic_vector(13 downto 0);
		sin    : out std_logic_vector(13 downto 0);
		cos    : out std_logic_vector(13 downto 0)
		);
end entity;

architecture rtl of sincos_lut_14 is

	signal pdsADD, pdcADD :  std_logic;
	signal dsADD, dcADD :  std_logic;
	signal sAz, cAz   :  std_logic;
	signal sADD, cADD :  std_logic_vector(13 DOWNTO 0);
	signal msin, mcos :  std_logic_vector(13 DOWNTO 0);

	type rom_mem is array (0 to 4095) of std_logic_vector (15 downto 0);
	constant isin : rom_mem :=(  
    x"0000", x"0003", x"0006", x"0009", x"000d", x"0010", x"0013", x"0016", 
    x"0019", x"001c", x"001f", x"0023", x"0026", x"0029", x"002c", x"002f", 
    x"0032", x"0035", x"0039", x"003c", x"003f", x"0042", x"0045", x"0048", 
    x"004b", x"004f", x"0052", x"0055", x"0058", x"005b", x"005e", x"0061", 
    x"0065", x"0068", x"006b", x"006e", x"0071", x"0074", x"0077", x"007b", 
    x"007e", x"0081", x"0084", x"0087", x"008a", x"008d", x"0090", x"0094", 
    x"0097", x"009a", x"009d", x"00a0", x"00a3", x"00a6", x"00aa", x"00ad", 
    x"00b0", x"00b3", x"00b6", x"00b9", x"00bc", x"00c0", x"00c3", x"00c6", 
    x"00c9", x"00cc", x"00cf", x"00d2", x"00d6", x"00d9", x"00dc", x"00df", 
    x"00e2", x"00e5", x"00e8", x"00ec", x"00ef", x"00f2", x"00f5", x"00f8", 
    x"00fb", x"00fe", x"0102", x"0105", x"0108", x"010b", x"010e", x"0111", 
    x"0114", x"0118", x"011b", x"011e", x"0121", x"0124", x"0127", x"012a", 
    x"012d", x"0131", x"0134", x"0137", x"013a", x"013d", x"0140", x"0143", 
    x"0147", x"014a", x"014d", x"0150", x"0153", x"0156", x"0159", x"015d", 
    x"0160", x"0163", x"0166", x"0169", x"016c", x"016f", x"0173", x"0176", 
    x"0179", x"017c", x"017f", x"0182", x"0185", x"0189", x"018c", x"018f", 
    x"0192", x"0195", x"0198", x"019b", x"019e", x"01a2", x"01a5", x"01a8", 
    x"01ab", x"01ae", x"01b1", x"01b4", x"01b8", x"01bb", x"01be", x"01c1", 
    x"01c4", x"01c7", x"01ca", x"01ce", x"01d1", x"01d4", x"01d7", x"01da", 
    x"01dd", x"01e0", x"01e3", x"01e7", x"01ea", x"01ed", x"01f0", x"01f3", 
    x"01f6", x"01f9", x"01fd", x"0200", x"0203", x"0206", x"0209", x"020c", 
    x"020f", x"0212", x"0216", x"0219", x"021c", x"021f", x"0222", x"0225", 
    x"0228", x"022c", x"022f", x"0232", x"0235", x"0238", x"023b", x"023e", 
    x"0242", x"0245", x"0248", x"024b", x"024e", x"0251", x"0254", x"0257", 
    x"025b", x"025e", x"0261", x"0264", x"0267", x"026a", x"026d", x"0270", 
    x"0274", x"0277", x"027a", x"027d", x"0280", x"0283", x"0286", x"028a", 
    x"028d", x"0290", x"0293", x"0296", x"0299", x"029c", x"029f", x"02a3", 
    x"02a6", x"02a9", x"02ac", x"02af", x"02b2", x"02b5", x"02b9", x"02bc", 
    x"02bf", x"02c2", x"02c5", x"02c8", x"02cb", x"02ce", x"02d2", x"02d5", 
    x"02d8", x"02db", x"02de", x"02e1", x"02e4", x"02e7", x"02eb", x"02ee", 
    x"02f1", x"02f4", x"02f7", x"02fa", x"02fd", x"0300", x"0304", x"0307", 
    x"030a", x"030d", x"0310", x"0313", x"0316", x"0319", x"031d", x"0320", 
    x"0323", x"0326", x"0329", x"032c", x"032f", x"0332", x"0336", x"0339", 
    x"033c", x"033f", x"0342", x"0345", x"0348", x"034b", x"034f", x"0352", 
    x"0355", x"0358", x"035b", x"035e", x"0361", x"0364", x"0368", x"036b", 
    x"036e", x"0371", x"0374", x"0377", x"037a", x"037d", x"0381", x"0384", 
    x"0387", x"038a", x"038d", x"0390", x"0393", x"0396", x"039a", x"039d", 
    x"03a0", x"03a3", x"03a6", x"03a9", x"03ac", x"03af", x"03b3", x"03b6", 
    x"03b9", x"03bc", x"03bf", x"03c2", x"03c5", x"03c8", x"03cb", x"03cf", 
    x"03d2", x"03d5", x"03d8", x"03db", x"03de", x"03e1", x"03e4", x"03e8", 
    x"03eb", x"03ee", x"03f1", x"03f4", x"03f7", x"03fa", x"03fd", x"0400", 
    x"0404", x"0407", x"040a", x"040d", x"0410", x"0413", x"0416", x"0419", 
    x"041d", x"0420", x"0423", x"0426", x"0429", x"042c", x"042f", x"0432", 
    x"0435", x"0439", x"043c", x"043f", x"0442", x"0445", x"0448", x"044b", 
    x"044e", x"0451", x"0455", x"0458", x"045b", x"045e", x"0461", x"0464", 
    x"0467", x"046a", x"046d", x"0471", x"0474", x"0477", x"047a", x"047d", 
    x"0480", x"0483", x"0486", x"0489", x"048d", x"0490", x"0493", x"0496", 
    x"0499", x"049c", x"049f", x"04a2", x"04a5", x"04a9", x"04ac", x"04af", 
    x"04b2", x"04b5", x"04b8", x"04bb", x"04be", x"04c1", x"04c5", x"04c8", 
    x"04cb", x"04ce", x"04d1", x"04d4", x"04d7", x"04da", x"04dd", x"04e0", 
    x"04e4", x"04e7", x"04ea", x"04ed", x"04f0", x"04f3", x"04f6", x"04f9", 
    x"04fc", x"04ff", x"0503", x"0506", x"0509", x"050c", x"050f", x"0512", 
    x"0515", x"0518", x"051b", x"051f", x"0522", x"0525", x"0528", x"052b", 
    x"052e", x"0531", x"0534", x"0537", x"053a", x"053e", x"0541", x"0544", 
    x"0547", x"054a", x"054d", x"0550", x"0553", x"0556", x"0559", x"055c", 
    x"0560", x"0563", x"0566", x"0569", x"056c", x"056f", x"0572", x"0575", 
    x"0578", x"057b", x"057f", x"0582", x"0585", x"0588", x"058b", x"058e", 
    x"0591", x"0594", x"0597", x"059a", x"059d", x"05a1", x"05a4", x"05a7", 
    x"05aa", x"05ad", x"05b0", x"05b3", x"05b6", x"05b9", x"05bc", x"05bf", 
    x"05c3", x"05c6", x"05c9", x"05cc", x"05cf", x"05d2", x"05d5", x"05d8", 
    x"05db", x"05de", x"05e1", x"05e5", x"05e8", x"05eb", x"05ee", x"05f1", 
    x"05f4", x"05f7", x"05fa", x"05fd", x"0600", x"0603", x"0606", x"060a", 
    x"060d", x"0610", x"0613", x"0616", x"0619", x"061c", x"061f", x"0622", 
    x"0625", x"0628", x"062b", x"062f", x"0632", x"0635", x"0638", x"063b", 
    x"063e", x"0641", x"0644", x"0647", x"064a", x"064d", x"0650", x"0654", 
    x"0657", x"065a", x"065d", x"0660", x"0663", x"0666", x"0669", x"066c", 
    x"066f", x"0672", x"0675", x"0678", x"067c", x"067f", x"0682", x"0685", 
    x"0688", x"068b", x"068e", x"0691", x"0694", x"0697", x"069a", x"069d", 
    x"06a0", x"06a4", x"06a7", x"06aa", x"06ad", x"06b0", x"06b3", x"06b6", 
    x"06b9", x"06bc", x"06bf", x"06c2", x"06c5", x"06c8", x"06cb", x"06cf", 
    x"06d2", x"06d5", x"06d8", x"06db", x"06de", x"06e1", x"06e4", x"06e7", 
    x"06ea", x"06ed", x"06f0", x"06f3", x"06f6", x"06f9", x"06fd", x"0700", 
    x"0703", x"0706", x"0709", x"070c", x"070f", x"0712", x"0715", x"0718", 
    x"071b", x"071e", x"0721", x"0724", x"0727", x"072a", x"072e", x"0731", 
    x"0734", x"0737", x"073a", x"073d", x"0740", x"0743", x"0746", x"0749", 
    x"074c", x"074f", x"0752", x"0755", x"0758", x"075b", x"075e", x"0762", 
    x"0765", x"0768", x"076b", x"076e", x"0771", x"0774", x"0777", x"077a", 
    x"077d", x"0780", x"0783", x"0786", x"0789", x"078c", x"078f", x"0792", 
    x"0795", x"0799", x"079c", x"079f", x"07a2", x"07a5", x"07a8", x"07ab", 
    x"07ae", x"07b1", x"07b4", x"07b7", x"07ba", x"07bd", x"07c0", x"07c3", 
    x"07c6", x"07c9", x"07cc", x"07cf", x"07d2", x"07d5", x"07d9", x"07dc", 
    x"07df", x"07e2", x"07e5", x"07e8", x"07eb", x"07ee", x"07f1", x"07f4", 
    x"07f7", x"07fa", x"07fd", x"0800", x"0803", x"0806", x"0809", x"080c", 
    x"080f", x"0812", x"0815", x"0818", x"081b", x"081e", x"0822", x"0825", 
    x"0828", x"082b", x"082e", x"0831", x"0834", x"0837", x"083a", x"083d", 
    x"0840", x"0843", x"0846", x"0849", x"084c", x"084f", x"0852", x"0855", 
    x"0858", x"085b", x"085e", x"0861", x"0864", x"0867", x"086a", x"086d", 
    x"0870", x"0873", x"0876", x"087a", x"087d", x"0880", x"0883", x"0886", 
    x"0889", x"088c", x"088f", x"0892", x"0895", x"0898", x"089b", x"089e", 
    x"08a1", x"08a4", x"08a7", x"08aa", x"08ad", x"08b0", x"08b3", x"08b6", 
    x"08b9", x"08bc", x"08bf", x"08c2", x"08c5", x"08c8", x"08cb", x"08ce", 
    x"08d1", x"08d4", x"08d7", x"08da", x"08dd", x"08e0", x"08e3", x"08e6", 
    x"08e9", x"08ec", x"08ef", x"08f2", x"08f5", x"08f8", x"08fb", x"08fe", 
    x"0901", x"0904", x"0908", x"090b", x"090e", x"0911", x"0914", x"0917", 
    x"091a", x"091d", x"0920", x"0923", x"0926", x"0929", x"092c", x"092f", 
    x"0932", x"0935", x"0938", x"093b", x"093e", x"0941", x"0944", x"0947", 
    x"094a", x"094d", x"0950", x"0953", x"0956", x"0959", x"095c", x"095f", 
    x"0962", x"0965", x"0968", x"096b", x"096e", x"0971", x"0974", x"0977", 
    x"097a", x"097d", x"0980", x"0983", x"0986", x"0989", x"098c", x"098f", 
    x"0992", x"0995", x"0998", x"099b", x"099e", x"09a1", x"09a4", x"09a7", 
    x"09aa", x"09ad", x"09b0", x"09b3", x"09b6", x"09b9", x"09bc", x"09bf", 
    x"09c2", x"09c5", x"09c8", x"09cb", x"09ce", x"09d1", x"09d4", x"09d7", 
    x"09da", x"09dd", x"09e0", x"09e3", x"09e6", x"09e9", x"09ec", x"09ef", 
    x"09f1", x"09f4", x"09f7", x"09fa", x"09fd", x"0a00", x"0a03", x"0a06", 
    x"0a09", x"0a0c", x"0a0f", x"0a12", x"0a15", x"0a18", x"0a1b", x"0a1e", 
    x"0a21", x"0a24", x"0a27", x"0a2a", x"0a2d", x"0a30", x"0a33", x"0a36", 
    x"0a39", x"0a3c", x"0a3f", x"0a42", x"0a45", x"0a48", x"0a4b", x"0a4e", 
    x"0a51", x"0a54", x"0a57", x"0a5a", x"0a5d", x"0a60", x"0a63", x"0a66", 
    x"0a69", x"0a6c", x"0a6f", x"0a72", x"0a74", x"0a77", x"0a7a", x"0a7d", 
    x"0a80", x"0a83", x"0a86", x"0a89", x"0a8c", x"0a8f", x"0a92", x"0a95", 
    x"0a98", x"0a9b", x"0a9e", x"0aa1", x"0aa4", x"0aa7", x"0aaa", x"0aad", 
    x"0ab0", x"0ab3", x"0ab6", x"0ab9", x"0abc", x"0abf", x"0ac2", x"0ac5", 
    x"0ac7", x"0aca", x"0acd", x"0ad0", x"0ad3", x"0ad6", x"0ad9", x"0adc", 
    x"0adf", x"0ae2", x"0ae5", x"0ae8", x"0aeb", x"0aee", x"0af1", x"0af4", 
    x"0af7", x"0afa", x"0afd", x"0b00", x"0b03", x"0b05", x"0b08", x"0b0b", 
    x"0b0e", x"0b11", x"0b14", x"0b17", x"0b1a", x"0b1d", x"0b20", x"0b23", 
    x"0b26", x"0b29", x"0b2c", x"0b2f", x"0b32", x"0b35", x"0b38", x"0b3a", 
    x"0b3d", x"0b40", x"0b43", x"0b46", x"0b49", x"0b4c", x"0b4f", x"0b52", 
    x"0b55", x"0b58", x"0b5b", x"0b5e", x"0b61", x"0b64", x"0b67", x"0b6a", 
    x"0b6c", x"0b6f", x"0b72", x"0b75", x"0b78", x"0b7b", x"0b7e", x"0b81", 
    x"0b84", x"0b87", x"0b8a", x"0b8d", x"0b90", x"0b93", x"0b95", x"0b98", 
    x"0b9b", x"0b9e", x"0ba1", x"0ba4", x"0ba7", x"0baa", x"0bad", x"0bb0", 
    x"0bb3", x"0bb6", x"0bb9", x"0bbc", x"0bbe", x"0bc1", x"0bc4", x"0bc7", 
    x"0bca", x"0bcd", x"0bd0", x"0bd3", x"0bd6", x"0bd9", x"0bdc", x"0bdf", 
    x"0be1", x"0be4", x"0be7", x"0bea", x"0bed", x"0bf0", x"0bf3", x"0bf6", 
    x"0bf9", x"0bfc", x"0bff", x"0c02", x"0c04", x"0c07", x"0c0a", x"0c0d", 
    x"0c10", x"0c13", x"0c16", x"0c19", x"0c1c", x"0c1f", x"0c22", x"0c24", 
    x"0c27", x"0c2a", x"0c2d", x"0c30", x"0c33", x"0c36", x"0c39", x"0c3c", 
    x"0c3f", x"0c41", x"0c44", x"0c47", x"0c4a", x"0c4d", x"0c50", x"0c53", 
    x"0c56", x"0c59", x"0c5c", x"0c5e", x"0c61", x"0c64", x"0c67", x"0c6a", 
    x"0c6d", x"0c70", x"0c73", x"0c76", x"0c79", x"0c7b", x"0c7e", x"0c81", 
    x"0c84", x"0c87", x"0c8a", x"0c8d", x"0c90", x"0c93", x"0c95", x"0c98", 
    x"0c9b", x"0c9e", x"0ca1", x"0ca4", x"0ca7", x"0caa", x"0cad", x"0caf", 
    x"0cb2", x"0cb5", x"0cb8", x"0cbb", x"0cbe", x"0cc1", x"0cc4", x"0cc6", 
    x"0cc9", x"0ccc", x"0ccf", x"0cd2", x"0cd5", x"0cd8", x"0cdb", x"0cdd", 
    x"0ce0", x"0ce3", x"0ce6", x"0ce9", x"0cec", x"0cef", x"0cf2", x"0cf4", 
    x"0cf7", x"0cfa", x"0cfd", x"0d00", x"0d03", x"0d06", x"0d09", x"0d0b", 
    x"0d0e", x"0d11", x"0d14", x"0d17", x"0d1a", x"0d1d", x"0d1f", x"0d22", 
    x"0d25", x"0d28", x"0d2b", x"0d2e", x"0d31", x"0d34", x"0d36", x"0d39", 
    x"0d3c", x"0d3f", x"0d42", x"0d45", x"0d48", x"0d4a", x"0d4d", x"0d50", 
    x"0d53", x"0d56", x"0d59", x"0d5c", x"0d5e", x"0d61", x"0d64", x"0d67", 
    x"0d6a", x"0d6d", x"0d70", x"0d72", x"0d75", x"0d78", x"0d7b", x"0d7e", 
    x"0d81", x"0d83", x"0d86", x"0d89", x"0d8c", x"0d8f", x"0d92", x"0d95", 
    x"0d97", x"0d9a", x"0d9d", x"0da0", x"0da3", x"0da6", x"0da8", x"0dab", 
    x"0dae", x"0db1", x"0db4", x"0db7", x"0db9", x"0dbc", x"0dbf", x"0dc2", 
    x"0dc5", x"0dc8", x"0dca", x"0dcd", x"0dd0", x"0dd3", x"0dd6", x"0dd9", 
    x"0ddb", x"0dde", x"0de1", x"0de4", x"0de7", x"0dea", x"0dec", x"0def", 
    x"0df2", x"0df5", x"0df8", x"0dfb", x"0dfd", x"0e00", x"0e03", x"0e06", 
    x"0e09", x"0e0c", x"0e0e", x"0e11", x"0e14", x"0e17", x"0e1a", x"0e1c", 
    x"0e1f", x"0e22", x"0e25", x"0e28", x"0e2b", x"0e2d", x"0e30", x"0e33", 
    x"0e36", x"0e39", x"0e3b", x"0e3e", x"0e41", x"0e44", x"0e47", x"0e49", 
    x"0e4c", x"0e4f", x"0e52", x"0e55", x"0e58", x"0e5a", x"0e5d", x"0e60", 
    x"0e63", x"0e66", x"0e68", x"0e6b", x"0e6e", x"0e71", x"0e74", x"0e76", 
    x"0e79", x"0e7c", x"0e7f", x"0e82", x"0e84", x"0e87", x"0e8a", x"0e8d", 
    x"0e90", x"0e92", x"0e95", x"0e98", x"0e9b", x"0e9e", x"0ea0", x"0ea3", 
    x"0ea6", x"0ea9", x"0eac", x"0eae", x"0eb1", x"0eb4", x"0eb7", x"0eb9", 
    x"0ebc", x"0ebf", x"0ec2", x"0ec5", x"0ec7", x"0eca", x"0ecd", x"0ed0", 
    x"0ed3", x"0ed5", x"0ed8", x"0edb", x"0ede", x"0ee0", x"0ee3", x"0ee6", 
    x"0ee9", x"0eec", x"0eee", x"0ef1", x"0ef4", x"0ef7", x"0ef9", x"0efc", 
    x"0eff", x"0f02", x"0f05", x"0f07", x"0f0a", x"0f0d", x"0f10", x"0f12", 
    x"0f15", x"0f18", x"0f1b", x"0f1e", x"0f20", x"0f23", x"0f26", x"0f29", 
    x"0f2b", x"0f2e", x"0f31", x"0f34", x"0f36", x"0f39", x"0f3c", x"0f3f", 
    x"0f41", x"0f44", x"0f47", x"0f4a", x"0f4d", x"0f4f", x"0f52", x"0f55", 
    x"0f58", x"0f5a", x"0f5d", x"0f60", x"0f63", x"0f65", x"0f68", x"0f6b", 
    x"0f6e", x"0f70", x"0f73", x"0f76", x"0f79", x"0f7b", x"0f7e", x"0f81", 
    x"0f84", x"0f86", x"0f89", x"0f8c", x"0f8f", x"0f91", x"0f94", x"0f97", 
    x"0f9a", x"0f9c", x"0f9f", x"0fa2", x"0fa4", x"0fa7", x"0faa", x"0fad", 
    x"0faf", x"0fb2", x"0fb5", x"0fb8", x"0fba", x"0fbd", x"0fc0", x"0fc3", 
    x"0fc5", x"0fc8", x"0fcb", x"0fce", x"0fd0", x"0fd3", x"0fd6", x"0fd8", 
    x"0fdb", x"0fde", x"0fe1", x"0fe3", x"0fe6", x"0fe9", x"0fec", x"0fee", 
    x"0ff1", x"0ff4", x"0ff6", x"0ff9", x"0ffc", x"0fff", x"1001", x"1004", 
    x"1007", x"1009", x"100c", x"100f", x"1012", x"1014", x"1017", x"101a", 
    x"101c", x"101f", x"1022", x"1025", x"1027", x"102a", x"102d", x"102f", 
    x"1032", x"1035", x"1038", x"103a", x"103d", x"1040", x"1042", x"1045", 
    x"1048", x"104b", x"104d", x"1050", x"1053", x"1055", x"1058", x"105b", 
    x"105d", x"1060", x"1063", x"1066", x"1068", x"106b", x"106e", x"1070", 
    x"1073", x"1076", x"1078", x"107b", x"107e", x"1080", x"1083", x"1086", 
    x"1089", x"108b", x"108e", x"1091", x"1093", x"1096", x"1099", x"109b", 
    x"109e", x"10a1", x"10a3", x"10a6", x"10a9", x"10ab", x"10ae", x"10b1", 
    x"10b3", x"10b6", x"10b9", x"10bc", x"10be", x"10c1", x"10c4", x"10c6", 
    x"10c9", x"10cc", x"10ce", x"10d1", x"10d4", x"10d6", x"10d9", x"10dc", 
    x"10de", x"10e1", x"10e4", x"10e6", x"10e9", x"10ec", x"10ee", x"10f1", 
    x"10f4", x"10f6", x"10f9", x"10fc", x"10fe", x"1101", x"1104", x"1106", 
    x"1109", x"110c", x"110e", x"1111", x"1114", x"1116", x"1119", x"111c", 
    x"111e", x"1121", x"1123", x"1126", x"1129", x"112b", x"112e", x"1131", 
    x"1133", x"1136", x"1139", x"113b", x"113e", x"1141", x"1143", x"1146", 
    x"1149", x"114b", x"114e", x"1150", x"1153", x"1156", x"1158", x"115b", 
    x"115e", x"1160", x"1163", x"1166", x"1168", x"116b", x"116d", x"1170", 
    x"1173", x"1175", x"1178", x"117b", x"117d", x"1180", x"1183", x"1185", 
    x"1188", x"118a", x"118d", x"1190", x"1192", x"1195", x"1198", x"119a", 
    x"119d", x"119f", x"11a2", x"11a5", x"11a7", x"11aa", x"11ad", x"11af", 
    x"11b2", x"11b4", x"11b7", x"11ba", x"11bc", x"11bf", x"11c1", x"11c4", 
    x"11c7", x"11c9", x"11cc", x"11cf", x"11d1", x"11d4", x"11d6", x"11d9", 
    x"11dc", x"11de", x"11e1", x"11e3", x"11e6", x"11e9", x"11eb", x"11ee", 
    x"11f0", x"11f3", x"11f6", x"11f8", x"11fb", x"11fd", x"1200", x"1203", 
    x"1205", x"1208", x"120a", x"120d", x"1210", x"1212", x"1215", x"1217", 
    x"121a", x"121c", x"121f", x"1222", x"1224", x"1227", x"1229", x"122c", 
    x"122f", x"1231", x"1234", x"1236", x"1239", x"123c", x"123e", x"1241", 
    x"1243", x"1246", x"1248", x"124b", x"124e", x"1250", x"1253", x"1255", 
    x"1258", x"125a", x"125d", x"1260", x"1262", x"1265", x"1267", x"126a", 
    x"126c", x"126f", x"1272", x"1274", x"1277", x"1279", x"127c", x"127e", 
    x"1281", x"1284", x"1286", x"1289", x"128b", x"128e", x"1290", x"1293", 
    x"1295", x"1298", x"129b", x"129d", x"12a0", x"12a2", x"12a5", x"12a7", 
    x"12aa", x"12ac", x"12af", x"12b2", x"12b4", x"12b7", x"12b9", x"12bc", 
    x"12be", x"12c1", x"12c3", x"12c6", x"12c8", x"12cb", x"12ce", x"12d0", 
    x"12d3", x"12d5", x"12d8", x"12da", x"12dd", x"12df", x"12e2", x"12e4", 
    x"12e7", x"12e9", x"12ec", x"12ef", x"12f1", x"12f4", x"12f6", x"12f9", 
    x"12fb", x"12fe", x"1300", x"1303", x"1305", x"1308", x"130a", x"130d", 
    x"130f", x"1312", x"1314", x"1317", x"1319", x"131c", x"131e", x"1321", 
    x"1324", x"1326", x"1329", x"132b", x"132e", x"1330", x"1333", x"1335", 
    x"1338", x"133a", x"133d", x"133f", x"1342", x"1344", x"1347", x"1349", 
    x"134c", x"134e", x"1351", x"1353", x"1356", x"1358", x"135b", x"135d", 
    x"1360", x"1362", x"1365", x"1367", x"136a", x"136c", x"136f", x"1371", 
    x"1374", x"1376", x"1379", x"137b", x"137e", x"1380", x"1383", x"1385", 
    x"1388", x"138a", x"138d", x"138f", x"1392", x"1394", x"1397", x"1399", 
    x"139c", x"139e", x"13a0", x"13a3", x"13a5", x"13a8", x"13aa", x"13ad", 
    x"13af", x"13b2", x"13b4", x"13b7", x"13b9", x"13bc", x"13be", x"13c1", 
    x"13c3", x"13c6", x"13c8", x"13cb", x"13cd", x"13cf", x"13d2", x"13d4", 
    x"13d7", x"13d9", x"13dc", x"13de", x"13e1", x"13e3", x"13e6", x"13e8", 
    x"13eb", x"13ed", x"13ef", x"13f2", x"13f4", x"13f7", x"13f9", x"13fc", 
    x"13fe", x"1401", x"1403", x"1406", x"1408", x"140a", x"140d", x"140f", 
    x"1412", x"1414", x"1417", x"1419", x"141c", x"141e", x"1420", x"1423", 
    x"1425", x"1428", x"142a", x"142d", x"142f", x"1432", x"1434", x"1436", 
    x"1439", x"143b", x"143e", x"1440", x"1443", x"1445", x"1447", x"144a", 
    x"144c", x"144f", x"1451", x"1454", x"1456", x"1458", x"145b", x"145d", 
    x"1460", x"1462", x"1465", x"1467", x"1469", x"146c", x"146e", x"1471", 
    x"1473", x"1475", x"1478", x"147a", x"147d", x"147f", x"1482", x"1484", 
    x"1486", x"1489", x"148b", x"148e", x"1490", x"1492", x"1495", x"1497", 
    x"149a", x"149c", x"149e", x"14a1", x"14a3", x"14a6", x"14a8", x"14aa", 
    x"14ad", x"14af", x"14b2", x"14b4", x"14b6", x"14b9", x"14bb", x"14be", 
    x"14c0", x"14c2", x"14c5", x"14c7", x"14ca", x"14cc", x"14ce", x"14d1", 
    x"14d3", x"14d5", x"14d8", x"14da", x"14dd", x"14df", x"14e1", x"14e4", 
    x"14e6", x"14e9", x"14eb", x"14ed", x"14f0", x"14f2", x"14f4", x"14f7", 
    x"14f9", x"14fc", x"14fe", x"1500", x"1503", x"1505", x"1507", x"150a", 
    x"150c", x"150e", x"1511", x"1513", x"1516", x"1518", x"151a", x"151d", 
    x"151f", x"1521", x"1524", x"1526", x"1528", x"152b", x"152d", x"152f", 
    x"1532", x"1534", x"1537", x"1539", x"153b", x"153e", x"1540", x"1542", 
    x"1545", x"1547", x"1549", x"154c", x"154e", x"1550", x"1553", x"1555", 
    x"1557", x"155a", x"155c", x"155e", x"1561", x"1563", x"1565", x"1568", 
    x"156a", x"156c", x"156f", x"1571", x"1573", x"1576", x"1578", x"157a", 
    x"157d", x"157f", x"1581", x"1584", x"1586", x"1588", x"158b", x"158d", 
    x"158f", x"1592", x"1594", x"1596", x"1599", x"159b", x"159d", x"15a0", 
    x"15a2", x"15a4", x"15a7", x"15a9", x"15ab", x"15ad", x"15b0", x"15b2", 
    x"15b4", x"15b7", x"15b9", x"15bb", x"15be", x"15c0", x"15c2", x"15c5", 
    x"15c7", x"15c9", x"15cb", x"15ce", x"15d0", x"15d2", x"15d5", x"15d7", 
    x"15d9", x"15db", x"15de", x"15e0", x"15e2", x"15e5", x"15e7", x"15e9", 
    x"15ec", x"15ee", x"15f0", x"15f2", x"15f5", x"15f7", x"15f9", x"15fc", 
    x"15fe", x"1600", x"1602", x"1605", x"1607", x"1609", x"160b", x"160e", 
    x"1610", x"1612", x"1615", x"1617", x"1619", x"161b", x"161e", x"1620", 
    x"1622", x"1624", x"1627", x"1629", x"162b", x"162e", x"1630", x"1632", 
    x"1634", x"1637", x"1639", x"163b", x"163d", x"1640", x"1642", x"1644", 
    x"1646", x"1649", x"164b", x"164d", x"164f", x"1652", x"1654", x"1656", 
    x"1658", x"165b", x"165d", x"165f", x"1661", x"1664", x"1666", x"1668", 
    x"166a", x"166d", x"166f", x"1671", x"1673", x"1676", x"1678", x"167a", 
    x"167c", x"167e", x"1681", x"1683", x"1685", x"1687", x"168a", x"168c", 
    x"168e", x"1690", x"1693", x"1695", x"1697", x"1699", x"169b", x"169e", 
    x"16a0", x"16a2", x"16a4", x"16a7", x"16a9", x"16ab", x"16ad", x"16af", 
    x"16b2", x"16b4", x"16b6", x"16b8", x"16bb", x"16bd", x"16bf", x"16c1", 
    x"16c3", x"16c6", x"16c8", x"16ca", x"16cc", x"16ce", x"16d1", x"16d3", 
    x"16d5", x"16d7", x"16d9", x"16dc", x"16de", x"16e0", x"16e2", x"16e4", 
    x"16e7", x"16e9", x"16eb", x"16ed", x"16ef", x"16f2", x"16f4", x"16f6", 
    x"16f8", x"16fa", x"16fc", x"16ff", x"1701", x"1703", x"1705", x"1707", 
    x"170a", x"170c", x"170e", x"1710", x"1712", x"1714", x"1717", x"1719", 
    x"171b", x"171d", x"171f", x"1721", x"1724", x"1726", x"1728", x"172a", 
    x"172c", x"172e", x"1731", x"1733", x"1735", x"1737", x"1739", x"173b", 
    x"173e", x"1740", x"1742", x"1744", x"1746", x"1748", x"174b", x"174d", 
    x"174f", x"1751", x"1753", x"1755", x"1757", x"175a", x"175c", x"175e", 
    x"1760", x"1762", x"1764", x"1766", x"1769", x"176b", x"176d", x"176f", 
    x"1771", x"1773", x"1775", x"1778", x"177a", x"177c", x"177e", x"1780", 
    x"1782", x"1784", x"1787", x"1789", x"178b", x"178d", x"178f", x"1791", 
    x"1793", x"1795", x"1798", x"179a", x"179c", x"179e", x"17a0", x"17a2", 
    x"17a4", x"17a6", x"17a8", x"17ab", x"17ad", x"17af", x"17b1", x"17b3", 
    x"17b5", x"17b7", x"17b9", x"17bb", x"17be", x"17c0", x"17c2", x"17c4", 
    x"17c6", x"17c8", x"17ca", x"17cc", x"17ce", x"17d0", x"17d3", x"17d5", 
    x"17d7", x"17d9", x"17db", x"17dd", x"17df", x"17e1", x"17e3", x"17e5", 
    x"17e8", x"17ea", x"17ec", x"17ee", x"17f0", x"17f2", x"17f4", x"17f6", 
    x"17f8", x"17fa", x"17fc", x"17fe", x"1800", x"1803", x"1805", x"1807", 
    x"1809", x"180b", x"180d", x"180f", x"1811", x"1813", x"1815", x"1817", 
    x"1819", x"181b", x"181d", x"1820", x"1822", x"1824", x"1826", x"1828", 
    x"182a", x"182c", x"182e", x"1830", x"1832", x"1834", x"1836", x"1838", 
    x"183a", x"183c", x"183e", x"1840", x"1842", x"1845", x"1847", x"1849", 
    x"184b", x"184d", x"184f", x"1851", x"1853", x"1855", x"1857", x"1859", 
    x"185b", x"185d", x"185f", x"1861", x"1863", x"1865", x"1867", x"1869", 
    x"186b", x"186d", x"186f", x"1871", x"1873", x"1875", x"1877", x"1879", 
    x"187b", x"187e", x"1880", x"1882", x"1884", x"1886", x"1888", x"188a", 
    x"188c", x"188e", x"1890", x"1892", x"1894", x"1896", x"1898", x"189a", 
    x"189c", x"189e", x"18a0", x"18a2", x"18a4", x"18a6", x"18a8", x"18aa", 
    x"18ac", x"18ae", x"18b0", x"18b2", x"18b4", x"18b6", x"18b8", x"18ba", 
    x"18bc", x"18be", x"18c0", x"18c2", x"18c4", x"18c6", x"18c8", x"18ca", 
    x"18cc", x"18ce", x"18d0", x"18d2", x"18d4", x"18d6", x"18d8", x"18da", 
    x"18db", x"18dd", x"18df", x"18e1", x"18e3", x"18e5", x"18e7", x"18e9", 
    x"18eb", x"18ed", x"18ef", x"18f1", x"18f3", x"18f5", x"18f7", x"18f9", 
    x"18fb", x"18fd", x"18ff", x"1901", x"1903", x"1905", x"1907", x"1909", 
    x"190b", x"190d", x"190f", x"1911", x"1913", x"1914", x"1916", x"1918", 
    x"191a", x"191c", x"191e", x"1920", x"1922", x"1924", x"1926", x"1928", 
    x"192a", x"192c", x"192e", x"1930", x"1932", x"1934", x"1935", x"1937", 
    x"1939", x"193b", x"193d", x"193f", x"1941", x"1943", x"1945", x"1947", 
    x"1949", x"194b", x"194d", x"194f", x"1950", x"1952", x"1954", x"1956", 
    x"1958", x"195a", x"195c", x"195e", x"1960", x"1962", x"1964", x"1966", 
    x"1967", x"1969", x"196b", x"196d", x"196f", x"1971", x"1973", x"1975", 
    x"1977", x"1979", x"197b", x"197c", x"197e", x"1980", x"1982", x"1984", 
    x"1986", x"1988", x"198a", x"198c", x"198d", x"198f", x"1991", x"1993", 
    x"1995", x"1997", x"1999", x"199b", x"199d", x"199e", x"19a0", x"19a2", 
    x"19a4", x"19a6", x"19a8", x"19aa", x"19ac", x"19ad", x"19af", x"19b1", 
    x"19b3", x"19b5", x"19b7", x"19b9", x"19bb", x"19bc", x"19be", x"19c0", 
    x"19c2", x"19c4", x"19c6", x"19c8", x"19c9", x"19cb", x"19cd", x"19cf", 
    x"19d1", x"19d3", x"19d5", x"19d6", x"19d8", x"19da", x"19dc", x"19de", 
    x"19e0", x"19e2", x"19e3", x"19e5", x"19e7", x"19e9", x"19eb", x"19ed", 
    x"19ee", x"19f0", x"19f2", x"19f4", x"19f6", x"19f8", x"19f9", x"19fb", 
    x"19fd", x"19ff", x"1a01", x"1a03", x"1a04", x"1a06", x"1a08", x"1a0a", 
    x"1a0c", x"1a0e", x"1a0f", x"1a11", x"1a13", x"1a15", x"1a17", x"1a19", 
    x"1a1a", x"1a1c", x"1a1e", x"1a20", x"1a22", x"1a23", x"1a25", x"1a27", 
    x"1a29", x"1a2b", x"1a2c", x"1a2e", x"1a30", x"1a32", x"1a34", x"1a35", 
    x"1a37", x"1a39", x"1a3b", x"1a3d", x"1a3e", x"1a40", x"1a42", x"1a44", 
    x"1a46", x"1a47", x"1a49", x"1a4b", x"1a4d", x"1a4f", x"1a50", x"1a52", 
    x"1a54", x"1a56", x"1a58", x"1a59", x"1a5b", x"1a5d", x"1a5f", x"1a60", 
    x"1a62", x"1a64", x"1a66", x"1a68", x"1a69", x"1a6b", x"1a6d", x"1a6f", 
    x"1a70", x"1a72", x"1a74", x"1a76", x"1a77", x"1a79", x"1a7b", x"1a7d", 
    x"1a7f", x"1a80", x"1a82", x"1a84", x"1a86", x"1a87", x"1a89", x"1a8b", 
    x"1a8d", x"1a8e", x"1a90", x"1a92", x"1a94", x"1a95", x"1a97", x"1a99", 
    x"1a9b", x"1a9c", x"1a9e", x"1aa0", x"1aa2", x"1aa3", x"1aa5", x"1aa7", 
    x"1aa8", x"1aaa", x"1aac", x"1aae", x"1aaf", x"1ab1", x"1ab3", x"1ab5", 
    x"1ab6", x"1ab8", x"1aba", x"1abc", x"1abd", x"1abf", x"1ac1", x"1ac2", 
    x"1ac4", x"1ac6", x"1ac8", x"1ac9", x"1acb", x"1acd", x"1ace", x"1ad0", 
    x"1ad2", x"1ad4", x"1ad5", x"1ad7", x"1ad9", x"1ada", x"1adc", x"1ade", 
    x"1ae0", x"1ae1", x"1ae3", x"1ae5", x"1ae6", x"1ae8", x"1aea", x"1aeb", 
    x"1aed", x"1aef", x"1af1", x"1af2", x"1af4", x"1af6", x"1af7", x"1af9", 
    x"1afb", x"1afc", x"1afe", x"1b00", x"1b01", x"1b03", x"1b05", x"1b07", 
    x"1b08", x"1b0a", x"1b0c", x"1b0d", x"1b0f", x"1b11", x"1b12", x"1b14", 
    x"1b16", x"1b17", x"1b19", x"1b1b", x"1b1c", x"1b1e", x"1b20", x"1b21", 
    x"1b23", x"1b25", x"1b26", x"1b28", x"1b2a", x"1b2b", x"1b2d", x"1b2f", 
    x"1b30", x"1b32", x"1b34", x"1b35", x"1b37", x"1b39", x"1b3a", x"1b3c", 
    x"1b3d", x"1b3f", x"1b41", x"1b42", x"1b44", x"1b46", x"1b47", x"1b49", 
    x"1b4b", x"1b4c", x"1b4e", x"1b50", x"1b51", x"1b53", x"1b54", x"1b56", 
    x"1b58", x"1b59", x"1b5b", x"1b5d", x"1b5e", x"1b60", x"1b61", x"1b63", 
    x"1b65", x"1b66", x"1b68", x"1b6a", x"1b6b", x"1b6d", x"1b6e", x"1b70", 
    x"1b72", x"1b73", x"1b75", x"1b76", x"1b78", x"1b7a", x"1b7b", x"1b7d", 
    x"1b7f", x"1b80", x"1b82", x"1b83", x"1b85", x"1b87", x"1b88", x"1b8a", 
    x"1b8b", x"1b8d", x"1b8f", x"1b90", x"1b92", x"1b93", x"1b95", x"1b97", 
    x"1b98", x"1b9a", x"1b9b", x"1b9d", x"1b9e", x"1ba0", x"1ba2", x"1ba3", 
    x"1ba5", x"1ba6", x"1ba8", x"1baa", x"1bab", x"1bad", x"1bae", x"1bb0", 
    x"1bb1", x"1bb3", x"1bb5", x"1bb6", x"1bb8", x"1bb9", x"1bbb", x"1bbc", 
    x"1bbe", x"1bc0", x"1bc1", x"1bc3", x"1bc4", x"1bc6", x"1bc7", x"1bc9", 
    x"1bca", x"1bcc", x"1bce", x"1bcf", x"1bd1", x"1bd2", x"1bd4", x"1bd5", 
    x"1bd7", x"1bd8", x"1bda", x"1bdc", x"1bdd", x"1bdf", x"1be0", x"1be2", 
    x"1be3", x"1be5", x"1be6", x"1be8", x"1be9", x"1beb", x"1bec", x"1bee", 
    x"1bf0", x"1bf1", x"1bf3", x"1bf4", x"1bf6", x"1bf7", x"1bf9", x"1bfa", 
    x"1bfc", x"1bfd", x"1bff", x"1c00", x"1c02", x"1c03", x"1c05", x"1c06", 
    x"1c08", x"1c09", x"1c0b", x"1c0c", x"1c0e", x"1c0f", x"1c11", x"1c12", 
    x"1c14", x"1c15", x"1c17", x"1c18", x"1c1a", x"1c1b", x"1c1d", x"1c1e", 
    x"1c20", x"1c21", x"1c23", x"1c24", x"1c26", x"1c27", x"1c29", x"1c2a", 
    x"1c2c", x"1c2d", x"1c2f", x"1c30", x"1c32", x"1c33", x"1c35", x"1c36", 
    x"1c38", x"1c39", x"1c3b", x"1c3c", x"1c3e", x"1c3f", x"1c41", x"1c42", 
    x"1c44", x"1c45", x"1c47", x"1c48", x"1c4a", x"1c4b", x"1c4c", x"1c4e", 
    x"1c4f", x"1c51", x"1c52", x"1c54", x"1c55", x"1c57", x"1c58", x"1c5a", 
    x"1c5b", x"1c5d", x"1c5e", x"1c5f", x"1c61", x"1c62", x"1c64", x"1c65", 
    x"1c67", x"1c68", x"1c6a", x"1c6b", x"1c6c", x"1c6e", x"1c6f", x"1c71", 
    x"1c72", x"1c74", x"1c75", x"1c77", x"1c78", x"1c79", x"1c7b", x"1c7c", 
    x"1c7e", x"1c7f", x"1c81", x"1c82", x"1c83", x"1c85", x"1c86", x"1c88", 
    x"1c89", x"1c8a", x"1c8c", x"1c8d", x"1c8f", x"1c90", x"1c92", x"1c93", 
    x"1c94", x"1c96", x"1c97", x"1c99", x"1c9a", x"1c9b", x"1c9d", x"1c9e", 
    x"1ca0", x"1ca1", x"1ca2", x"1ca4", x"1ca5", x"1ca7", x"1ca8", x"1ca9", 
    x"1cab", x"1cac", x"1cae", x"1caf", x"1cb0", x"1cb2", x"1cb3", x"1cb5", 
    x"1cb6", x"1cb7", x"1cb9", x"1cba", x"1cbc", x"1cbd", x"1cbe", x"1cc0", 
    x"1cc1", x"1cc2", x"1cc4", x"1cc5", x"1cc7", x"1cc8", x"1cc9", x"1ccb", 
    x"1ccc", x"1ccd", x"1ccf", x"1cd0", x"1cd1", x"1cd3", x"1cd4", x"1cd6", 
    x"1cd7", x"1cd8", x"1cda", x"1cdb", x"1cdc", x"1cde", x"1cdf", x"1ce0", 
    x"1ce2", x"1ce3", x"1ce4", x"1ce6", x"1ce7", x"1ce9", x"1cea", x"1ceb", 
    x"1ced", x"1cee", x"1cef", x"1cf1", x"1cf2", x"1cf3", x"1cf5", x"1cf6", 
    x"1cf7", x"1cf9", x"1cfa", x"1cfb", x"1cfd", x"1cfe", x"1cff", x"1d01", 
    x"1d02", x"1d03", x"1d05", x"1d06", x"1d07", x"1d09", x"1d0a", x"1d0b", 
    x"1d0c", x"1d0e", x"1d0f", x"1d10", x"1d12", x"1d13", x"1d14", x"1d16", 
    x"1d17", x"1d18", x"1d1a", x"1d1b", x"1d1c", x"1d1e", x"1d1f", x"1d20", 
    x"1d21", x"1d23", x"1d24", x"1d25", x"1d27", x"1d28", x"1d29", x"1d2a", 
    x"1d2c", x"1d2d", x"1d2e", x"1d30", x"1d31", x"1d32", x"1d34", x"1d35", 
    x"1d36", x"1d37", x"1d39", x"1d3a", x"1d3b", x"1d3c", x"1d3e", x"1d3f", 
    x"1d40", x"1d42", x"1d43", x"1d44", x"1d45", x"1d47", x"1d48", x"1d49", 
    x"1d4a", x"1d4c", x"1d4d", x"1d4e", x"1d4f", x"1d51", x"1d52", x"1d53", 
    x"1d55", x"1d56", x"1d57", x"1d58", x"1d5a", x"1d5b", x"1d5c", x"1d5d", 
    x"1d5f", x"1d60", x"1d61", x"1d62", x"1d64", x"1d65", x"1d66", x"1d67", 
    x"1d68", x"1d6a", x"1d6b", x"1d6c", x"1d6d", x"1d6f", x"1d70", x"1d71", 
    x"1d72", x"1d74", x"1d75", x"1d76", x"1d77", x"1d78", x"1d7a", x"1d7b", 
    x"1d7c", x"1d7d", x"1d7f", x"1d80", x"1d81", x"1d82", x"1d83", x"1d85", 
    x"1d86", x"1d87", x"1d88", x"1d89", x"1d8b", x"1d8c", x"1d8d", x"1d8e", 
    x"1d8f", x"1d91", x"1d92", x"1d93", x"1d94", x"1d95", x"1d97", x"1d98", 
    x"1d99", x"1d9a", x"1d9b", x"1d9d", x"1d9e", x"1d9f", x"1da0", x"1da1", 
    x"1da3", x"1da4", x"1da5", x"1da6", x"1da7", x"1da8", x"1daa", x"1dab", 
    x"1dac", x"1dad", x"1dae", x"1db0", x"1db1", x"1db2", x"1db3", x"1db4", 
    x"1db5", x"1db7", x"1db8", x"1db9", x"1dba", x"1dbb", x"1dbc", x"1dbe", 
    x"1dbf", x"1dc0", x"1dc1", x"1dc2", x"1dc3", x"1dc4", x"1dc6", x"1dc7", 
    x"1dc8", x"1dc9", x"1dca", x"1dcb", x"1dcc", x"1dce", x"1dcf", x"1dd0", 
    x"1dd1", x"1dd2", x"1dd3", x"1dd4", x"1dd6", x"1dd7", x"1dd8", x"1dd9", 
    x"1dda", x"1ddb", x"1ddc", x"1dde", x"1ddf", x"1de0", x"1de1", x"1de2", 
    x"1de3", x"1de4", x"1de5", x"1de7", x"1de8", x"1de9", x"1dea", x"1deb", 
    x"1dec", x"1ded", x"1dee", x"1def", x"1df1", x"1df2", x"1df3", x"1df4", 
    x"1df5", x"1df6", x"1df7", x"1df8", x"1df9", x"1dfa", x"1dfc", x"1dfd", 
    x"1dfe", x"1dff", x"1e00", x"1e01", x"1e02", x"1e03", x"1e04", x"1e05", 
    x"1e06", x"1e08", x"1e09", x"1e0a", x"1e0b", x"1e0c", x"1e0d", x"1e0e", 
    x"1e0f", x"1e10", x"1e11", x"1e12", x"1e13", x"1e14", x"1e16", x"1e17", 
    x"1e18", x"1e19", x"1e1a", x"1e1b", x"1e1c", x"1e1d", x"1e1e", x"1e1f", 
    x"1e20", x"1e21", x"1e22", x"1e23", x"1e24", x"1e25", x"1e27", x"1e28", 
    x"1e29", x"1e2a", x"1e2b", x"1e2c", x"1e2d", x"1e2e", x"1e2f", x"1e30", 
    x"1e31", x"1e32", x"1e33", x"1e34", x"1e35", x"1e36", x"1e37", x"1e38", 
    x"1e39", x"1e3a", x"1e3b", x"1e3c", x"1e3d", x"1e3e", x"1e3f", x"1e40", 
    x"1e41", x"1e42", x"1e44", x"1e45", x"1e46", x"1e47", x"1e48", x"1e49", 
    x"1e4a", x"1e4b", x"1e4c", x"1e4d", x"1e4e", x"1e4f", x"1e50", x"1e51", 
    x"1e52", x"1e53", x"1e54", x"1e55", x"1e56", x"1e57", x"1e58", x"1e59", 
    x"1e5a", x"1e5b", x"1e5c", x"1e5d", x"1e5e", x"1e5f", x"1e60", x"1e61", 
    x"1e62", x"1e63", x"1e64", x"1e65", x"1e66", x"1e66", x"1e67", x"1e68", 
    x"1e69", x"1e6a", x"1e6b", x"1e6c", x"1e6d", x"1e6e", x"1e6f", x"1e70", 
    x"1e71", x"1e72", x"1e73", x"1e74", x"1e75", x"1e76", x"1e77", x"1e78", 
    x"1e79", x"1e7a", x"1e7b", x"1e7c", x"1e7d", x"1e7e", x"1e7f", x"1e80", 
    x"1e81", x"1e81", x"1e82", x"1e83", x"1e84", x"1e85", x"1e86", x"1e87", 
    x"1e88", x"1e89", x"1e8a", x"1e8b", x"1e8c", x"1e8d", x"1e8e", x"1e8f", 
    x"1e90", x"1e90", x"1e91", x"1e92", x"1e93", x"1e94", x"1e95", x"1e96", 
    x"1e97", x"1e98", x"1e99", x"1e9a", x"1e9b", x"1e9c", x"1e9c", x"1e9d", 
    x"1e9e", x"1e9f", x"1ea0", x"1ea1", x"1ea2", x"1ea3", x"1ea4", x"1ea5", 
    x"1ea6", x"1ea6", x"1ea7", x"1ea8", x"1ea9", x"1eaa", x"1eab", x"1eac", 
    x"1ead", x"1eae", x"1eaf", x"1eaf", x"1eb0", x"1eb1", x"1eb2", x"1eb3", 
    x"1eb4", x"1eb5", x"1eb6", x"1eb6", x"1eb7", x"1eb8", x"1eb9", x"1eba", 
    x"1ebb", x"1ebc", x"1ebd", x"1ebe", x"1ebe", x"1ebf", x"1ec0", x"1ec1", 
    x"1ec2", x"1ec3", x"1ec4", x"1ec4", x"1ec5", x"1ec6", x"1ec7", x"1ec8", 
    x"1ec9", x"1eca", x"1eca", x"1ecb", x"1ecc", x"1ecd", x"1ece", x"1ecf", 
    x"1ed0", x"1ed0", x"1ed1", x"1ed2", x"1ed3", x"1ed4", x"1ed5", x"1ed5", 
    x"1ed6", x"1ed7", x"1ed8", x"1ed9", x"1eda", x"1eda", x"1edb", x"1edc", 
    x"1edd", x"1ede", x"1edf", x"1edf", x"1ee0", x"1ee1", x"1ee2", x"1ee3", 
    x"1ee4", x"1ee4", x"1ee5", x"1ee6", x"1ee7", x"1ee8", x"1ee8", x"1ee9", 
    x"1eea", x"1eeb", x"1eec", x"1eec", x"1eed", x"1eee", x"1eef", x"1ef0", 
    x"1ef1", x"1ef1", x"1ef2", x"1ef3", x"1ef4", x"1ef4", x"1ef5", x"1ef6", 
    x"1ef7", x"1ef8", x"1ef8", x"1ef9", x"1efa", x"1efb", x"1efc", x"1efc", 
    x"1efd", x"1efe", x"1eff", x"1f00", x"1f00", x"1f01", x"1f02", x"1f03", 
    x"1f03", x"1f04", x"1f05", x"1f06", x"1f06", x"1f07", x"1f08", x"1f09", 
    x"1f0a", x"1f0a", x"1f0b", x"1f0c", x"1f0d", x"1f0d", x"1f0e", x"1f0f", 
    x"1f10", x"1f10", x"1f11", x"1f12", x"1f13", x"1f13", x"1f14", x"1f15", 
    x"1f16", x"1f16", x"1f17", x"1f18", x"1f19", x"1f19", x"1f1a", x"1f1b", 
    x"1f1c", x"1f1c", x"1f1d", x"1f1e", x"1f1e", x"1f1f", x"1f20", x"1f21", 
    x"1f21", x"1f22", x"1f23", x"1f24", x"1f24", x"1f25", x"1f26", x"1f26", 
    x"1f27", x"1f28", x"1f29", x"1f29", x"1f2a", x"1f2b", x"1f2b", x"1f2c", 
    x"1f2d", x"1f2e", x"1f2e", x"1f2f", x"1f30", x"1f30", x"1f31", x"1f32", 
    x"1f32", x"1f33", x"1f34", x"1f35", x"1f35", x"1f36", x"1f37", x"1f37", 
    x"1f38", x"1f39", x"1f39", x"1f3a", x"1f3b", x"1f3b", x"1f3c", x"1f3d", 
    x"1f3d", x"1f3e", x"1f3f", x"1f3f", x"1f40", x"1f41", x"1f41", x"1f42", 
    x"1f43", x"1f44", x"1f44", x"1f45", x"1f46", x"1f46", x"1f47", x"1f47", 
    x"1f48", x"1f49", x"1f49", x"1f4a", x"1f4b", x"1f4b", x"1f4c", x"1f4d", 
    x"1f4d", x"1f4e", x"1f4f", x"1f4f", x"1f50", x"1f51", x"1f51", x"1f52", 
    x"1f53", x"1f53", x"1f54", x"1f54", x"1f55", x"1f56", x"1f56", x"1f57", 
    x"1f58", x"1f58", x"1f59", x"1f5a", x"1f5a", x"1f5b", x"1f5b", x"1f5c", 
    x"1f5d", x"1f5d", x"1f5e", x"1f5f", x"1f5f", x"1f60", x"1f60", x"1f61", 
    x"1f62", x"1f62", x"1f63", x"1f63", x"1f64", x"1f65", x"1f65", x"1f66", 
    x"1f66", x"1f67", x"1f68", x"1f68", x"1f69", x"1f69", x"1f6a", x"1f6b", 
    x"1f6b", x"1f6c", x"1f6c", x"1f6d", x"1f6e", x"1f6e", x"1f6f", x"1f6f", 
    x"1f70", x"1f71", x"1f71", x"1f72", x"1f72", x"1f73", x"1f73", x"1f74", 
    x"1f75", x"1f75", x"1f76", x"1f76", x"1f77", x"1f77", x"1f78", x"1f79", 
    x"1f79", x"1f7a", x"1f7a", x"1f7b", x"1f7b", x"1f7c", x"1f7d", x"1f7d", 
    x"1f7e", x"1f7e", x"1f7f", x"1f7f", x"1f80", x"1f80", x"1f81", x"1f82", 
    x"1f82", x"1f83", x"1f83", x"1f84", x"1f84", x"1f85", x"1f85", x"1f86", 
    x"1f86", x"1f87", x"1f87", x"1f88", x"1f89", x"1f89", x"1f8a", x"1f8a", 
    x"1f8b", x"1f8b", x"1f8c", x"1f8c", x"1f8d", x"1f8d", x"1f8e", x"1f8e", 
    x"1f8f", x"1f8f", x"1f90", x"1f90", x"1f91", x"1f91", x"1f92", x"1f92", 
    x"1f93", x"1f93", x"1f94", x"1f94", x"1f95", x"1f95", x"1f96", x"1f96", 
    x"1f97", x"1f97", x"1f98", x"1f98", x"1f99", x"1f99", x"1f9a", x"1f9a", 
    x"1f9b", x"1f9b", x"1f9c", x"1f9c", x"1f9d", x"1f9d", x"1f9e", x"1f9e", 
    x"1f9f", x"1f9f", x"1fa0", x"1fa0", x"1fa1", x"1fa1", x"1fa2", x"1fa2", 
    x"1fa3", x"1fa3", x"1fa4", x"1fa4", x"1fa4", x"1fa5", x"1fa5", x"1fa6", 
    x"1fa6", x"1fa7", x"1fa7", x"1fa8", x"1fa8", x"1fa9", x"1fa9", x"1faa", 
    x"1faa", x"1faa", x"1fab", x"1fab", x"1fac", x"1fac", x"1fad", x"1fad", 
    x"1fae", x"1fae", x"1fae", x"1faf", x"1faf", x"1fb0", x"1fb0", x"1fb1", 
    x"1fb1", x"1fb1", x"1fb2", x"1fb2", x"1fb3", x"1fb3", x"1fb4", x"1fb4", 
    x"1fb4", x"1fb5", x"1fb5", x"1fb6", x"1fb6", x"1fb7", x"1fb7", x"1fb7", 
    x"1fb8", x"1fb8", x"1fb9", x"1fb9", x"1fb9", x"1fba", x"1fba", x"1fbb", 
    x"1fbb", x"1fbb", x"1fbc", x"1fbc", x"1fbd", x"1fbd", x"1fbd", x"1fbe", 
    x"1fbe", x"1fbf", x"1fbf", x"1fbf", x"1fc0", x"1fc0", x"1fc1", x"1fc1", 
    x"1fc1", x"1fc2", x"1fc2", x"1fc3", x"1fc3", x"1fc3", x"1fc4", x"1fc4", 
    x"1fc4", x"1fc5", x"1fc5", x"1fc6", x"1fc6", x"1fc6", x"1fc7", x"1fc7", 
    x"1fc7", x"1fc8", x"1fc8", x"1fc8", x"1fc9", x"1fc9", x"1fca", x"1fca", 
    x"1fca", x"1fcb", x"1fcb", x"1fcb", x"1fcc", x"1fcc", x"1fcc", x"1fcd", 
    x"1fcd", x"1fcd", x"1fce", x"1fce", x"1fce", x"1fcf", x"1fcf", x"1fcf", 
    x"1fd0", x"1fd0", x"1fd0", x"1fd1", x"1fd1", x"1fd1", x"1fd2", x"1fd2", 
    x"1fd2", x"1fd3", x"1fd3", x"1fd3", x"1fd4", x"1fd4", x"1fd4", x"1fd5", 
    x"1fd5", x"1fd5", x"1fd6", x"1fd6", x"1fd6", x"1fd7", x"1fd7", x"1fd7", 
    x"1fd8", x"1fd8", x"1fd8", x"1fd8", x"1fd9", x"1fd9", x"1fd9", x"1fda", 
    x"1fda", x"1fda", x"1fdb", x"1fdb", x"1fdb", x"1fdb", x"1fdc", x"1fdc", 
    x"1fdc", x"1fdd", x"1fdd", x"1fdd", x"1fdd", x"1fde", x"1fde", x"1fde", 
    x"1fdf", x"1fdf", x"1fdf", x"1fdf", x"1fe0", x"1fe0", x"1fe0", x"1fe1", 
    x"1fe1", x"1fe1", x"1fe1", x"1fe2", x"1fe2", x"1fe2", x"1fe2", x"1fe3", 
    x"1fe3", x"1fe3", x"1fe3", x"1fe4", x"1fe4", x"1fe4", x"1fe4", x"1fe5", 
    x"1fe5", x"1fe5", x"1fe5", x"1fe6", x"1fe6", x"1fe6", x"1fe6", x"1fe7", 
    x"1fe7", x"1fe7", x"1fe7", x"1fe8", x"1fe8", x"1fe8", x"1fe8", x"1fe9", 
    x"1fe9", x"1fe9", x"1fe9", x"1fe9", x"1fea", x"1fea", x"1fea", x"1fea", 
    x"1feb", x"1feb", x"1feb", x"1feb", x"1feb", x"1fec", x"1fec", x"1fec", 
    x"1fec", x"1fed", x"1fed", x"1fed", x"1fed", x"1fed", x"1fee", x"1fee", 
    x"1fee", x"1fee", x"1fee", x"1fef", x"1fef", x"1fef", x"1fef", x"1fef", 
    x"1ff0", x"1ff0", x"1ff0", x"1ff0", x"1ff0", x"1ff1", x"1ff1", x"1ff1", 
    x"1ff1", x"1ff1", x"1ff1", x"1ff2", x"1ff2", x"1ff2", x"1ff2", x"1ff2", 
    x"1ff3", x"1ff3", x"1ff3", x"1ff3", x"1ff3", x"1ff3", x"1ff4", x"1ff4", 
    x"1ff4", x"1ff4", x"1ff4", x"1ff4", x"1ff5", x"1ff5", x"1ff5", x"1ff5", 
    x"1ff5", x"1ff5", x"1ff5", x"1ff6", x"1ff6", x"1ff6", x"1ff6", x"1ff6", 
    x"1ff6", x"1ff6", x"1ff7", x"1ff7", x"1ff7", x"1ff7", x"1ff7", x"1ff7", 
    x"1ff7", x"1ff8", x"1ff8", x"1ff8", x"1ff8", x"1ff8", x"1ff8", x"1ff8", 
    x"1ff8", x"1ff9", x"1ff9", x"1ff9", x"1ff9", x"1ff9", x"1ff9", x"1ff9", 
    x"1ff9", x"1ffa", x"1ffa", x"1ffa", x"1ffa", x"1ffa", x"1ffa", x"1ffa", 
    x"1ffa", x"1ffa", x"1ffb", x"1ffb", x"1ffb", x"1ffb", x"1ffb", x"1ffb", 
    x"1ffb", x"1ffb", x"1ffb", x"1ffb", x"1ffc", x"1ffc", x"1ffc", x"1ffc", 
    x"1ffc", x"1ffc", x"1ffc", x"1ffc", x"1ffc", x"1ffc", x"1ffc", x"1ffc", 
    x"1ffd", x"1ffd", x"1ffd", x"1ffd", x"1ffd", x"1ffd", x"1ffd", x"1ffd", 
    x"1ffd", x"1ffd", x"1ffd", x"1ffd", x"1ffd", x"1ffd", x"1ffd", x"1ffe", 
    x"1ffe", x"1ffe", x"1ffe", x"1ffe", x"1ffe", x"1ffe", x"1ffe", x"1ffe", 
    x"1ffe", x"1ffe", x"1ffe", x"1ffe", x"1ffe", x"1ffe", x"1ffe", x"1ffe", 
    x"1ffe", x"1ffe", x"1ffe", x"1ffe", x"1fff", x"1fff", x"1fff", x"1fff", 
    x"1fff", x"1fff", x"1fff", x"1fff", x"1fff", x"1fff", x"1fff", x"1fff", 
    x"1fff", x"1fff", x"1fff", x"1fff", x"1fff", x"1fff", x"1fff", x"1fff", 
    x"1fff", x"1fff", x"1fff", x"1fff", x"1fff", x"1fff", x"1fff", x"1fff");

begin

process (clk_i)
BEGIN
	if (rising_edge (clk_i)) then
		dsADD <= pdsADD;
		dcADD <= pdcADD;
		if ((sADD = ("01" & x"000")) or (sADD = ("11" & x"000"))) then
			sAz <= '1';
		else
			sAz <= '0';
		end if;
		if ((cADD = ("00" & x"000")) or (cADD = ("10" & x"000"))) then
			cAz <= '1';
		else
			cAz <= '0';
		end if;
		if (addr_i(13 downto 12) = "00") then
			pdsADD <= '0';
			pdcADD <= '0';
			sADD <= "00" & addr_i(11 downto 0);
			cADD <= "00" & (x"0" - addr_i(11 downto 0));
		elsif (addr_i(13 downto 12) = "01") then
			pdsADD <= '0';
			pdcADD <= '1';
			sADD <= "01" & (x"0" - addr_i(11 downto 0));
			cADD <= "01" &  addr_i(11 downto 0);
		elsif (addr_i(13 downto 12) = "10") then
			pdsADD <= '1';
			pdcADD <= '1';
			sADD <= "10" & addr_i(11 downto 0);
			cADD <= "10" & (x"0" - addr_i(11 downto 0));
		else -- (addr_i(13 downto 12) = "11") then
			pdsADD <= '1';
			pdcADD <= '0';
			sADD <= "11" & (x"0" - addr_i(11 downto 0));
			cADD <= "11" & addr_i(11 downto 0);
		end if;
		msin <= isin(conv_integer(sADD(11 downto 0)))(13 downto 0);
		mcos <= isin(conv_integer(cADD(11 downto 0)))(13 downto 0);
		if (dsADD = '0') then
			if (sAz = '0') then
				sin <= msin(13 downto 0);
			else
				sin <= ("01" & x"fff");
			end if;
		else
			if (sAz = '0') then
				sin <= x"0" - msin(13 downto 0);
			else
				sin <= ("10" & x"001");
			end if;
			
		end if;
		if (dcADD = '0') then
			if (cAz = '0') then
				cos <= mcos(13 downto 0);
			else
				cos <= ("01" & x"fff");
			end if;			
		else 
			if (cAz = '0') then
				cos <= x"0" - mcos(13 downto 0);
			else
				cos <= ("10" & x"001");
			end if;
			
		end if;	
	end if;
end process;

end architecture;
